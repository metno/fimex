netcdf coordTest {
dimensions:
	time = UNLIMITED ; // (4 currently)
	sigma = 4 ;
	x = 11 ;
	y = 11 ;
variables:
	double time(time) ;
		time:long_name = "time" ;
		time:standard_name = "time" ;
		time:units = "seconds since 1970-01-01 00:00:00 +00:00" ;
	long forecast_reference_time ;
	    forecast_reference_time:standard_name = "forecast_reference_time" ;
		forecast_reference_time:units = "hours since 2000-01-01 00:00:00 +00:00" ;
	short sigma(sigma) ;
		sigma:description = "atmosphere sigma coordinate" ;
		sigma:long_name = "atmosphere_sigma_coordinate" ;
		sigma:standard_name = "atmosphere_sigma_coordinate" ;
		sigma:positive = "up" ;
		sigma:scale_factor = 0.001f ;
	int projection_1 ;
		projection_1:proj4 = "+proj=stere +lat_0=90 +lon_0=0 +lat_ts=60 +units=m +a=6.371e+06 +e=0 +no_defs" ;
		projection_1:grid_mapping_name = "stereographic" ;
		projection_1:scale_factor_at_projection_origin = 0.933012701907249 ;
		projection_1:longitude_of_projection_origin = 0. ;
		projection_1:latitude_of_projection_origin = 90. ;
	int x(x) ;
		x:long_name = "x-coordinate in Cartesian system" ;
		x:standard_name = "projection_x_coordinate" ;
		x:units = "m" ;
	int y(y) ;
		y:long_name = "y-coordinate in Cartesian system" ;
		y:standard_name = "projection_y_coordinate" ;
		y:units = "m" ;
	double longitude(y, x) ;
		longitude:units = "degree_east" ;
		longitude:long_name = "longitude" ;
		longitude:standard_name = "longitude" ;
	double latitude(y, x) ;
		latitude:units = "degree_north" ;
		latitude:long_name = "latitude" ;
		latitude:standard_name = "latitude" ;
	short altitude(time, y, x) ;
		altitude:_FillValue = -32767s ;
		altitude:long_name = "altitude" ;
		altitude:standard_name = "altitude" ;
		altitude:units = "m" ;
		altitude:grid_mapping = "projection_1" ;
		altitude:coordinates = "longitude latitude" ;
	short sea_surface_temperature(time, y, x) ;
		sea_surface_temperature:long_name = "sea_surface_temperature" ;
		sea_surface_temperature:standard_name = "sea_surface_temperature" ;
		sea_surface_temperature:units = "K" ;
		sea_surface_temperature:grid_mapping = "projection_1" ;
		sea_surface_temperature:coordinates = "longitude latitude" ;
		sea_surface_temperature:scale_factor = 0.01f ;
	float precipitation_amount(time, y, x) ;
		precipitation_amount:_FillValue = -32767.f ;
		precipitation_amount:long_name = "precipitation_amount" ;
		precipitation_amount:standard_name = "precipitation_amount" ;
		precipitation_amount:units = "kg/m2" ;
		precipitation_amount:grid_mapping = "projection_1" ;
		precipitation_amount:coordinates = "longitude latitude" ;
	short land_ice_area_fraction(time, y, x) ;
		land_ice_area_fraction:long_name = "land_ice_area_fraction" ;
		land_ice_area_fraction:metno_name = "land_ice_area_fraction" ;
		land_ice_area_fraction:scale_factor = 0.0001f ;
		land_ice_area_fraction:units = "1" ;
		land_ice_area_fraction:grid_mapping = "projection_1" ;
		land_ice_area_fraction:coordinates = "longitude latitude" ;
	short cloud_area_fraction(time, y, x) ;
		cloud_area_fraction:scale_factor = 0.0001f ;
		cloud_area_fraction:_FillValue = -32767s ;
		cloud_area_fraction:cell_methods = "time: point" ;
		cloud_area_fraction:long_name = "cloud_area_fraction" ;
		cloud_area_fraction:standard_name = "cloud_area_fraction" ;
		cloud_area_fraction:units = "1" ;
		cloud_area_fraction:grid_mapping = "projection_1" ;
		cloud_area_fraction:coordinates = "longitude latitude" ;
	short air_temperature(time, y, x) ;
		air_temperature:_FillValue = -32767s ;
		air_temperature:cell_methods = "time: point height: p" ;
		air_temperature:long_name = "air_temperature" ;
		air_temperature:standard_name = "air_temperature" ;
		air_temperature:units = "K" ;
		air_temperature:grid_mapping = "projection_1" ;
		air_temperature:coordinates = "longitude latitude" ;
		air_temperature:scale_factor = 0.01f ;
	float x_wind_10m(time, y, x) ;
		x_wind_10m:_FillValue = 9.96921e+36f ;
		x_wind_10m:cell_methods = "time: point height: 10m" ;
		x_wind_10m:long_name = "x_wind_10m" ;
		x_wind_10m:metno_name = "x_wind_10m" ;
		x_wind_10m:units = "m s-1" ;
		x_wind_10m:grid_mapping = "projection_1" ;
		x_wind_10m:coordinates = "longitude latitude" ;
	float y_wind_10m(time, y, x) ;
		y_wind_10m:_FillValue = 9.96921e+36f ;
		y_wind_10m:cell_methods = "time: point height: 10m" ;
		y_wind_10m:long_name = "y_wind_10m" ;
		y_wind_10m:standard_name = "y_wind_10m" ;
		y_wind_10m:units = "m s-1" ;
		y_wind_10m:grid_mapping = "projection_1" ;
		y_wind_10m:coordinates = "longitude latitude" ;
	short cloud_area_fraction_in_atmosphere_layer(time, sigma, y, x) ;
		cloud_area_fraction_in_atmosphere_layer:_FillValue = -32767s ;
		cloud_area_fraction_in_atmosphere_layer:long_name = "cloud_area_fraction_in_atmosphere_layer" ;
		cloud_area_fraction_in_atmosphere_layer:standard_name = "cloud_area_fraction_in_atmosphere_layer" ;
		cloud_area_fraction_in_atmosphere_layer:scale_factor = 0.0001f ;
		cloud_area_fraction_in_atmosphere_layer:units = "1" ;
		cloud_area_fraction_in_atmosphere_layer:grid_mapping = "projection_1" ;
		cloud_area_fraction_in_atmosphere_layer:coordinates = "longitude latitude" ;
	short sea_level_pressure(time, y, x) ;
		sea_level_pressure:scale_factor = 10.f ;
		sea_level_pressure:_FillValue = -32767s ;
		sea_level_pressure:cell_methods = "time: point" ;
		sea_level_pressure:long_name = "air_pressure_at_sea_level" ;
		sea_level_pressure:standard_name = "air_pressure_at_sea_level" ;
		sea_level_pressure:units = "Pa" ;
		sea_level_pressure:grid_mapping = "projection_1" ;
		sea_level_pressure:coordinates = "longitude latitude" ;
	short surface_snow_sickness(time, y, x) ;
		surface_snow_sickness:long_name = "surface_snow_sickness" ;
		surface_snow_sickness:standard_name = "surface_snow_sickness" ;
		surface_snow_sickness:units = "m" ;
		surface_snow_sickness:grid_mapping = "projection_1" ;
		surface_snow_sickness:coordinates = "longitude latitude" ;
		surface_snow_sickness:scale_factor = 0.001f ;

// global attributes:
		:Conventions = "CF-1.0" ;
		:institution = "Norwegian Meteorological Institute, met.no" ;
		:source = "HIRLAM" ;
		:title = "unknown" ;
		:min_time = "2007-05-16 00:00:00Z" ;
		:max_time = "2007-05-18" ;
		:Expires = "2007-06-15" ;
		:references = "unknown" ;
		:comment = "none" ;
		:history = "2010-02-09 creation by fimex from file \'../test/flth00.dat\'" ;
data:

 forecast_reference_time = 10 ;

 time = 1179309600, 1179313200, 1179316800, 1179320400 ;

 sigma = 300, 500, 850, 1000 ;

 projection_1 = _ ;

 x = -1705516, -1655353, -1605191, -1555029, -1504867, -1454704, -1404542, 
    -1354380, -1304218, -1254056, -1203893 ;

 y = -6872225, -6822063, -6771901, -6721738, -6671576, -6621414, -6571252, 
    -6521089, -6470927, -6420765, -6370603 ;

 longitude =
  -13.9377996159233, -13.5431788713008, -13.1472444238949, -12.7500277028342, 
    -12.3515608341056, -11.9518746349313, -11.5510085768871, 
    -11.1489928305179, -10.7458581694264, -10.341648062544, -9.93639050434804,
  -14.0362454440677, -13.6390538603117, -13.2405215536026, -12.8406804797004, 
    -12.4395633144029, -12.0372014343367, -11.6336349468322, 
    -11.2288946139368, -10.8230118219768, -10.4160307567415, -10.0079800409987,
  -14.1360633304441, -13.736269680603, -13.3351075574881, -12.932609453459, 
    -12.5288086050022, -12.1237369597633, -11.7174352740378, 
    -11.309934914639, -10.9012678947548, -10.4914791331451, -10.0805978964134,
  -14.2372825575012, -13.8348550758348, -13.4310306158913, -13.0258422167524, 
    -12.6193236866648, -12.2115075561413, -11.8024352439396, 
    -11.3921387352165, -10.9806506845137, -10.5680167600937, -10.1542668883725,
  -14.3399301378325, -13.9348365895563, -13.528316778696, -13.1204043013113, 
    -12.7111335486568, -12.3005376461761, -11.8886586888566, 
    -11.4755292940766, -11.0611827725664, -10.6456655590283, -10.2290082560918,
  -14.4440379376002, -14.0362455039508, -13.6269967173443, -13.2163257412266, 
    -12.8042675613046, -12.3908559102557, -11.9761335733649, 
    -11.5601338144382, -11.1428906156054, -10.7244511953915, -10.3048468495026,
  -14.5496345161434, -14.1391098919679, -13.7270979917868, -13.313633556964, 
    -12.8987521792745, -12.4824882111473, -12.0648851425071, 
    -11.645976898103, -11.2257981470302, -10.8043969094444, -10.3818051914367,
  -14.6567534563539, -14.2434627323742, -13.8286529477599, -13.4123594324664, 
    -12.9946183961435, -12.5754648237283, -12.1549429244323, 
    -11.7330872988008, -11.3099333188498, -10.8855298246393, -10.4599095504404,
  -14.7654249711455, -14.3493337340358, -13.9316907613006, -13.5125319822722, 
    -13.0918942364449, -12.6698131542321, -12.246333679056, 
    -11.8214911024267, -11.3953215156049, -10.9678745972713, -10.5391838281412,
  -14.8756844762093, -14.4567576880041, -14.0362455675766, -13.6141846545486, 
    -13.1906124304116, -12.7655651842582, -12.3390886089525, 
    -11.9112187024836, -11.4819922920831, -11.0514599142552, -10.6196558149333,
  -14.987563953486, -14.5657660542701, -14.1423482734753, -13.7173477720209, 
    -13.2908026856991, -12.8627499756907, -12.4332360998103, 
    -12.0022977783607, -11.5699725916495, -11.1363119536692, -10.7013508948374 ;

 latitude =
  28.4443934391326, 28.529204665858, 28.6116926308595, 28.6918393575517, 
    28.7696272800954, 28.8450396251899, 28.9180585743488, 28.9886686284868, 
    29.0568546497592, 29.1225999417882, 29.1858909572803,
  28.7913367354885, 28.8770436364891, 28.9604049318737, 29.0414022788004, 
    29.1200177516902, 29.1962342283441, 29.2700335328496, 29.3413998363176, 
    29.4103176781451, 29.4767700258027, 29.5407430332539,
  29.1393763014149, 29.2259910754273, 29.3102376524725, 29.3920973141981, 
    29.4715517661265, 29.5485835281654, 29.6231740578853, 29.6953071879173, 
    29.7649671263634, 29.8321364958657, 29.896801143551,
  29.4885110905519, 29.5760461637802, 29.661190198345, 29.7439240908398, 
    29.8242291684395, 29.9020875838766, 29.9774804188227, 30.050391158469, 
    30.120803670805, 30.1887002246833, 30.2540663520281,
  29.8387293862042, 29.92719738995, 30.0132512607874, 30.0968715004235, 
    30.1780390479492, 30.2567356793514, 30.3329420907311, 30.4066414105958, 
    30.4778171577228, 30.5464512379301, 30.6125288592987,
  30.1900331831424, 30.2794469961199, 30.366423326277, 30.4509422702881, 
    30.5329843691081, 30.6125310120951, 30.6895624997904, 30.7640615944649, 
    30.8360114562774, 30.9053936184553, 30.9721929562993,
  30.5424102551619, 30.6327829715716, 30.720694597394, 30.8061248138134, 
    30.8890537532864, 30.9694624083494, 31.0473306736818, 31.1226409354587, 
    31.1953759855087, 31.2655169746059, 31.3330484360362,
  30.8958621622374, 30.98720713544, 31.0760671493151, 31.1624214587625, 
    31.2462497770385, 31.3275326893276, 31.4062496738042, 31.4823827303536, 
    31.5559142724325, 31.6268250581628, 31.6950992692593,
  31.2503761456127, 31.3427069555009, 31.4325286741871, 31.5198201191576, 
    31.6045605734325, 31.6867302039798, 31.7663080614875, 31.8432757490271, 
    31.9176152913105, 31.9893070432765, 32.0583348251916,
  31.6059533058617, 31.6992838039532, 31.7900808127287, 31.8783227007689, 
    31.9639883094566, 32.0470573763152, 32.127508513197, 32.2053229154744, 
    32.2804822083842, 32.3529663327885, 32.422758737279,
  31.9625803272211, 32.0569246033144, 32.1487107236181, 32.2379165959552, 
    32.32452060831, 32.4085020571722, 32.489839103844, 32.5685125247556, 
    32.6445035345814, 32.7177916488523, 32.7883599339107 ;

 altitude =
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _ ;

 sea_surface_temperature =
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _ ;

 precipitation_amount =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0.001, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0.007, 0.008, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0.019, 0.009, 0.005, 0.001, 0, 0, 0, 0, 0, 0, 0,
  0.029, 0.014, 0.01, 0.001, 0, 0, 0, 0, 0, 0, 0,
  0.031, 0.028, 0.011, 0.001, 0, 0, 0, 0, 0, 0, 0,
  0.027, 0.038, 0.016, 0.007, 0.001, 0, 0, 0, 0, 0, 0,
  0.023, 0.033, 0.036, 0.017, 0.006, 0.001, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0.01, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0.02, 0.01, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0.03, 0.02, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0.04, 0.03, 0.02, 0, 0, 0, 0, 0, 0, 0, 0,
  0.04, 0.05, 0.03, 0.02, 0, 0, 0, 0, 0, 0, 0,
  0.03, 0.04, 0.04, 0.02, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0.01, 0.01, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0.03, 0.01, 0.01, 0, 0, 0, 0, 0, 0, 0, 0,
  0.04, 0.02, 0.01, 0, 0, 0, 0, 0, 0, 0, 0,
  0.05, 0.04, 0.01, 0, 0, 0, 0, 0, 0, 0, 0,
  0.03, 0.05, 0.02, 0.01, 0, 0, 0, 0, 0, 0, 0,
  0.03, 0.05, 0.04, 0.02, 0.01, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0.01, 0.01, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0.03, 0.01, 0.01, 0, 0, 0, 0, 0, 0, 0, 0,
  0.04, 0.02, 0.01, 0, 0, 0, 0, 0, 0, 0, 0,
  0.05, 0.04, 0.01, 0, 0, 0, 0, 0, 0, 0, 0,
  0.05, 0.05, 0.02, 0.01, 0, 0, 0, 0, 0, 0, 0,
  0.04, 0.05, 0.04, 0.02, 0.01, 0, 0, 0, 0, 0, 0 ;

 land_ice_area_fraction =
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _ ;

 cloud_area_fraction =
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 54, 157, 610, 552, 681,
  0, 0, 203, 78, 0, 297, 705, 569, 790, 717, 722,
  534, 698, 412, 80, 215, 893, 1108, 552, 526, 682, 436,
  150, 265, 410, 272, 556, 955, 806, 255, 153, 416, 82,
  692, 543, 1441, 1145, 912, 533, 103, 0, 4, 22, 1,
  7421, 7911, 6446, 3621, 2308, 2001, 1018, 0, 0, 0, 0,
  9684, 8305, 5208, 3730, 2692, 2102, 1047, 0, 0, 0, 0,
  6750, 4574, 2479, 2689, 1847, 932, 351, 0, 0, 0, 0,
  2126, 2867, 3740, 2226, 506, 0, 28, 0, 0, 0, 0,
  2905, 4522, 1367, 549, 81, 0, 0, 0, 0, 0, 0,
  4469, 5366, 1956, 45, 0, 0, 0, 0, 0, 0, 0,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _ ;

 air_temperature =
  29302, 29267, 29269, 29276, 29277, 29278, 29268, 29240, 29209, 29168, 29498,
  29264, 29297, 29275, 29277, 29282, 29280, 29269, 29248, 29222, 29181, 29390,
  29270, 29288, 29283, 29285, 29289, 29288, 29277, 29256, 29231, 29203, 29239,
  29274, 29273, 29285, 29289, 29292, 29294, 29285, 29262, 29237, 29223, 29175,
  29254, 29261, 29270, 29279, 29284, 29289, 29284, 29264, 29241, 29231, 29270,
  29218, 29221, 29232, 29246, 29254, 29264, 29266, 29253, 29232, 29210, 29236,
  29199, 29200, 29210, 29224, 29237, 29251, 29259, 29254, 29238, 29213, 29204,
  29191, 29192, 29200, 29213, 29230, 29248, 29261, 29265, 29259, 29243, 29220,
  29181, 29180, 29189, 29202, 29221, 29240, 29257, 29272, 29277, 29265, 29253,
  29172, 29168, 29175, 29191, 29208, 29228, 29249, 29271, 29285, 29282, 29275,
  29161, 29158, 29163, 29177, 29194, 29213, 29235, 29259, 29281, 29293, 29290,
  29337, 29280, 29275, 29281, 29282, 29283, 29274, 29244, 29207, 29185, 29618,
  29280, 29330, 29290, 29282, 29286, 29285, 29274, 29252, 29225, 29186, 29461,
  29281, 29309, 29294, 29293, 29296, 29294, 29283, 29261, 29235, 29207, 29264,
  29286, 29282, 29293, 29300, 29302, 29303, 29293, 29267, 29240, 29231, 29174,
  29269, 29272, 29281, 29291, 29296, 29300, 29293, 29267, 29241, 29239, 29269,
  29231, 29235, 29245, 29257, 29267, 29277, 29275, 29257, 29232, 29216, 29254,
  29208, 29213, 29226, 29239, 29252, 29264, 29269, 29260, 29240, 29217, 29223,
  29196, 29203, 29216, 29230, 29245, 29261, 29272, 29273, 29263, 29244, 29222,
  29187, 29191, 29200, 29216, 29232, 29252, 29271, 29282, 29280, 29266, 29255,
  29177, 29180, 29188, 29202, 29221, 29240, 29264, 29285, 29292, 29286, 29279,
  29170, 29170, 29177, 29191, 29207, 29227, 29251, 29276, 29294, 29298, 29294,
  29364, 29292, 29282, 29292, 29291, 29290, 29280, 29246, 29208, 29206, 29741,
  29288, 29355, 29300, 29289, 29294, 29292, 29280, 29255, 29225, 29189, 29533,
  29287, 29326, 29306, 29300, 29303, 29302, 29287, 29261, 29237, 29205, 29286,
  29294, 29291, 29305, 29307, 29310, 29311, 29296, 29267, 29245, 29235, 29170,
  29278, 29285, 29292, 29298, 29304, 29308, 29299, 29273, 29247, 29248, 29275,
  29238, 29247, 29257, 29268, 29280, 29285, 29281, 29264, 29237, 29226, 29276,
  29217, 29226, 29234, 29248, 29264, 29275, 29276, 29265, 29243, 29223, 29244,
  29208, 29216, 29225, 29238, 29257, 29274, 29282, 29278, 29263, 29244, 29231,
  29200, 29204, 29218, 29232, 29248, 29267, 29283, 29289, 29281, 29268, 29258,
  29191, 29193, 29208, 29222, 29235, 29256, 29279, 29293, 29295, 29287, 29280,
  29179, 29182, 29193, 29207, 29221, 29242, 29265, 29286, 29300, 29298, 29295,
  29380, 29302, 29289, 29294, 29295, 29293, 29281, 29248, 29212, 29209, 29765,
  29294, 29371, 29309, 29296, 29299, 29295, 29283, 29258, 29229, 29195, 29543,
  29293, 29337, 29312, 29306, 29308, 29305, 29290, 29265, 29241, 29213, 29293,
  29303, 29298, 29310, 29312, 29314, 29313, 29298, 29271, 29249, 29243, 29175,
  29289, 29293, 29299, 29303, 29309, 29311, 29300, 29274, 29250, 29252, 29263,
  29249, 29257, 29265, 29274, 29285, 29290, 29283, 29263, 29239, 29229, 29269,
  29228, 29236, 29244, 29257, 29271, 29281, 29278, 29263, 29243, 29226, 29247,
  29222, 29227, 29235, 29249, 29266, 29282, 29285, 29276, 29262, 29249, 29239,
  29215, 29218, 29226, 29239, 29258, 29278, 29289, 29288, 29281, 29271, 29267,
  29201, 29207, 29217, 29229, 29247, 29267, 29284, 29293, 29294, 29289, 29288,
  29187, 29195, 29205, 29216, 29231, 29251, 29272, 29290, 29300, 29300, 29300 ;

 x_wind_10m =
  -3.357, -2.556, -1.83, -1.413, -1.304, -1.311, -1.326, -1.16, -0.339, 
    1.146, 2.047,
  -3.615, -2.673, -2.006, -1.652, -1.673, -1.803, -1.921, -1.939, -1.191, 
    1.052, 2.539,
  -4.066, -3.291, -2.6, -2.317, -2.404, -2.632, -2.865, -3.017, -2.615, 
    -0.781, 1.471,
  -4.647, -4.059, -3.449, -3.221, -3.316, -3.581, -3.863, -4.094, -4.106, 
    -3.173, -0.3,
  -5.28, -4.757, -4.335, -4.12, -4.187, -4.428, -4.695, -4.979, -5.197, 
    -4.66, -1.721,
  -5.903, -5.393, -4.989, -4.79, -4.776, -5.034, -5.402, -5.751, -6.136, 
    -6.262, -5,
  -6.408, -5.887, -5.526, -5.286, -5.314, -5.577, -5.991, -6.469, -6.971, 
    -7.433, -7.47,
  -6.718, -6.269, -6.039, -5.743, -5.786, -5.992, -6.435, -7.092, -7.659, 
    -8.057, -8.252,
  -6.88, -6.612, -6.581, -6.278, -6.135, -6.201, -6.703, -7.499, -8.105, 
    -8.383, -8.121,
  -7.172, -7.007, -7.063, -6.825, -6.539, -6.43, -6.762, -7.5, -8.238, 
    -8.592, -8.424,
  -7.605, -7.368, -7.336, -7.345, -7.121, -6.884, -6.885, -7.251, -7.906, 
    -8.552, -8.83,
  -3.121, -2.288, -1.684, -1.386, -1.213, -1.085, -1.008, -0.727, 0.24, 1.66, 
    2.529,
  -3.248, -2.41, -1.862, -1.654, -1.584, -1.536, -1.555, -1.49, -0.663, 
    1.581, 3.083,
  -3.69, -3.013, -2.434, -2.267, -2.293, -2.356, -2.491, -2.585, -2.048, 
    -0.153, 2.105,
  -4.295, -3.81, -3.242, -3.09, -3.158, -3.29, -3.481, -3.648, -3.459, 
    -2.406, 0.449,
  -4.937, -4.562, -4.083, -3.938, -3.971, -4.116, -4.306, -4.483, -4.506, 
    -3.796, -0.881,
  -5.543, -5.159, -4.736, -4.602, -4.537, -4.815, -5.212, -5.368, -5.43, 
    -5.463, -4.38,
  -5.962, -5.642, -5.197, -5.06, -5.126, -5.508, -5.937, -6.167, -6.396, 
    -6.788, -7.061,
  -6.357, -5.983, -5.583, -5.408, -5.684, -6.084, -6.428, -6.814, -7.26, 
    -7.555, -7.905,
  -6.823, -6.227, -6.036, -5.802, -6.075, -6.389, -6.73, -7.26, -7.776, 
    -7.951, -7.723,
  -7.137, -6.657, -6.604, -6.45, -6.379, -6.383, -6.795, -7.557, -8.156, 
    -8.313, -7.872,
  -7.457, -7.1, -7.126, -7.067, -6.775, -6.518, -6.752, -7.488, -8.251, 
    -8.599, -8.352,
  -2.886, -2.015, -1.535, -1.369, -1.135, -0.864, -0.682, -0.317, 0.691, 
    2.169, 3.003,
  -2.887, -2.12, -1.713, -1.658, -1.497, -1.276, -1.199, -1.053, -0.156, 
    2.137, 3.619,
  -3.305, -2.726, -2.262, -2.217, -2.164, -2.079, -2.135, -2.154, -1.493, 
    0.483, 2.739,
  -3.943, -3.479, -3.044, -2.948, -2.959, -2.993, -3.131, -3.239, -2.877, 
    -1.654, 1.19,
  -4.594, -4.147, -3.862, -3.7, -3.692, -3.787, -3.949, -4.089, -3.916, 
    -2.943, -0.051,
  -5.1, -4.709, -4.464, -4.266, -4.211, -4.485, -4.857, -4.962, -4.855, 
    -4.777, -3.479,
  -5.652, -5.286, -4.979, -4.749, -4.664, -5.118, -5.71, -5.889, -5.842, 
    -6.058, -6.126,
  -6.243, -5.904, -5.36, -5.093, -5.101, -5.706, -6.394, -6.682, -6.713, 
    -6.663, -7.077,
  -6.807, -6.497, -5.605, -5.294, -5.531, -6.221, -6.823, -7.108, -7.247, 
    -7.178, -7.229,
  -7.241, -6.834, -5.996, -5.667, -5.887, -6.444, -7.041, -7.528, -7.812, 
    -7.733, -7.502,
  -7.438, -7.061, -6.524, -6.182, -6.201, -6.486, -7.061, -7.776, -8.261, 
    -8.285, -8.005,
  -2.494, -1.702, -1.277, -1.089, -0.877, -0.661, -0.505, -0.17, 0.727, 
    2.037, 2.994,
  -2.447, -1.796, -1.468, -1.373, -1.231, -1.066, -0.979, -0.797, -0.005, 
    1.929, 3.471,
  -2.871, -2.378, -2.008, -1.959, -1.93, -1.863, -1.86, -1.792, -1.16, 0.563, 
    2.706,
  -3.522, -3.11, -2.771, -2.712, -2.732, -2.72, -2.768, -2.807, -2.426, 
    -1.236, 1.364,
  -4.186, -3.785, -3.55, -3.433, -3.42, -3.407, -3.461, -3.61, -3.497, -2.48, 
    0.23,
  -4.744, -4.412, -4.034, -3.885, -3.928, -4.086, -4.248, -4.351, -4.385, 
    -4.155, -2.769,
  -5.2, -4.97, -4.674, -4.359, -4.347, -4.684, -5.055, -5.202, -5.249, 
    -5.409, -5.271,
  -5.665, -5.576, -5.331, -4.769, -4.696, -5.232, -5.851, -6.103, -6.063, 
    -6.11, -6.476,
  -6.212, -6.245, -5.753, -5.003, -5.019, -5.791, -6.586, -6.871, -6.753, 
    -6.672, -6.982,
  -6.744, -6.684, -5.928, -5.222, -5.51, -6.379, -7.127, -7.469, -7.484, 
    -7.332, -7.437,
  -7.028, -6.926, -6.258, -5.598, -5.92, -6.711, -7.424, -7.922, -8.178, 
    -8.106, -8.013 ;

 y_wind_10m =
  -8.136, -8.931, -9.331, -9.544, -9.757, -9.749, -9.4, -8.493, -6.057, 
    -1.274, -0.009,
  -8.426, -8.616, -9.407, -9.71, -9.973, -10.074, -9.837, -9.115, -6.835, 
    -1.896, 0.085,
  -8.612, -8.899, -9.566, -9.961, -10.301, -10.524, -10.508, -10.174, -8.76, 
    -4.804, -0.698,
  -8.856, -9.385, -9.87, -10.334, -10.747, -11.06, -11.183, -11.143, -10.71, 
    -8.539, -3.467,
  -9.16, -9.745, -10.243, -10.718, -11.193, -11.526, -11.617, -11.584, 
    -11.57, -11.096, -8.395,
  -9.382, -9.869, -10.343, -10.777, -11.237, -11.506, -11.629, -11.744, 
    -11.891, -12.132, -11.753,
  -9.338, -9.696, -10.186, -10.692, -11.01, -11.158, -11.218, -11.256, 
    -11.314, -11.469, -11.719,
  -9.179, -9.46, -10.004, -10.575, -10.806, -10.872, -10.764, -10.534, 
    -10.354, -10.073, -9.612,
  -9.073, -9.387, -9.954, -10.461, -10.846, -10.958, -10.728, -10.306, 
    -9.915, -9.509, -8.754,
  -9.022, -9.45, -9.709, -10.193, -10.644, -10.919, -10.946, -10.592, -9.872, 
    -9.12, -8.483,
  -8.921, -9.36, -9.485, -9.769, -10.151, -10.577, -10.891, -10.778, -10.058, 
    -9.069, -8.493,
  -8.079, -8.763, -9.167, -9.406, -9.5, -9.379, -9.014, -8.109, -5.812, 
    -1.524, -0.172,
  -8.3, -8.466, -9.207, -9.564, -9.703, -9.661, -9.4, -8.659, -6.481, -2.126, 
    -0.259,
  -8.446, -8.7, -9.301, -9.735, -10.011, -10.11, -10.046, -9.709, -8.326, 
    -4.759, -1.192,
  -8.663, -9.125, -9.592, -10.075, -10.454, -10.652, -10.73, -10.746, 
    -10.293, -8.192, -3.876,
  -8.953, -9.502, -10.057, -10.542, -10.926, -11.138, -11.227, -11.3, 
    -11.285, -10.715, -8.437,
  -9.193, -9.832, -10.354, -10.762, -11.074, -11.315, -11.46, -11.545, 
    -11.726, -12.019, -11.734,
  -9.167, -9.752, -10.253, -10.549, -10.791, -11.028, -11.15, -11.13, 
    -11.143, -11.393, -11.849,
  -9.08, -9.554, -10.039, -10.296, -10.514, -10.647, -10.604, -10.404, 
    -10.133, -9.869, -9.868,
  -9.11, -9.514, -9.977, -10.368, -10.648, -10.623, -10.34, -10.022, -9.762, 
    -9.403, -8.841,
  -9.101, -9.317, -9.692, -10.227, -10.575, -10.659, -10.413, -9.986, -9.613, 
    -9.221, -8.563,
  -8.933, -9.156, -9.411, -9.847, -10.239, -10.555, -10.565, -10.177, -9.606, 
    -9.076, -8.574,
  -8.01, -8.596, -8.997, -9.265, -9.239, -9.009, -8.633, -7.72, -5.562, 
    -1.782, -0.362,
  -8.165, -8.301, -8.99, -9.412, -9.42, -9.234, -8.957, -8.199, -6.127, 
    -2.343, -0.597,
  -8.25, -8.482, -9.027, -9.534, -9.709, -9.655, -9.555, -9.22, -7.887, 
    -4.694, -1.66,
  -8.477, -8.884, -9.341, -9.839, -10.15, -10.221, -10.244, -10.274, -9.809, 
    -7.852, -4.254,
  -8.843, -9.331, -9.92, -10.337, -10.664, -10.787, -10.813, -10.883, 
    -10.839, -10.374, -8.426,
  -9.15, -9.839, -10.324, -10.706, -10.964, -11.076, -11.141, -11.288, 
    -11.538, -11.768, -11.57,
  -9.125, -9.836, -10.352, -10.588, -10.724, -10.816, -10.885, -10.971, 
    -11.134, -11.437, -11.896,
  -9.04, -9.675, -10.178, -10.269, -10.332, -10.397, -10.4, -10.295, -10.15, 
    -10.17, -10.235,
  -9.111, -9.672, -10.013, -10.161, -10.298, -10.355, -10.249, -9.996, 
    -9.728, -9.563, -9.2,
  -8.987, -9.311, -9.789, -10.187, -10.394, -10.421, -10.195, -9.896, -9.716, 
    -9.447, -9.02,
  -8.886, -9.086, -9.506, -10.028, -10.404, -10.529, -10.315, -9.962, -9.674, 
    -9.322, -9.059,
  -8.154, -8.765, -9.128, -9.277, -9.222, -9.038, -8.681, -7.791, -5.766, 
    -2.171, -0.677,
  -8.277, -8.463, -9.145, -9.439, -9.42, -9.286, -9.028, -8.286, -6.321, 
    -2.712, -0.835,
  -8.372, -8.573, -9.162, -9.572, -9.712, -9.709, -9.609, -9.235, -8.001, 
    -5.029, -2.022,
  -8.594, -9, -9.442, -9.916, -10.179, -10.251, -10.25, -10.206, -9.806, 
    -8.11, -4.843,
  -8.943, -9.526, -9.992, -10.485, -10.767, -10.798, -10.791, -10.816, 
    -10.747, -10.509, -9.133,
  -9.25, -9.859, -10.383, -10.912, -11.187, -11.209, -11.226, -11.329, 
    -11.471, -11.845, -12.158,
  -9.16, -9.741, -10.434, -10.943, -11.071, -10.989, -10.989, -11.159, 
    -11.395, -11.742, -12.486,
  -9.026, -9.585, -10.311, -10.681, -10.645, -10.506, -10.485, -10.62, 
    -10.774, -10.776, -10.94,
  -9.135, -9.708, -10.214, -10.377, -10.359, -10.379, -10.415, -10.391, 
    -10.313, -10.145, -9.879,
  -9.131, -9.646, -10.065, -10.234, -10.428, -10.487, -10.425, -10.338, 
    -10.235, -10.06, -9.758,
  -9.108, -9.458, -9.886, -10.254, -10.577, -10.588, -10.383, -10.17, 
    -10.009, -9.883, -9.762 ;

 cloud_area_fraction_in_atmosphere_layer =
  0, 1, 2, 3, 4, 5, 6, 7, 8, 9, 10,
  11, 12, 13, 14, 15, 16, 17, 18, 19, 20, 21,
  22, 23, 24, 25, 26, 27, 28, 29, 30, 31, 32,
  33, 34, 35, 36, 37, 38, 39, 40, 41, 42, 43,
  44, 45, 46, 47, 48, 49, 50, 51, 52, 53, 54,
  55, 56, 57, 58, 59, 60, 61, 62, 63, 64, 65,
  66, 67, 68, 69, 70, 71, 72, 73, 74, 75, 76,
  77, 78, 79, 80, 81, 82, 83, 84, 85, 86, 87,
  88, 89, 90, 91, 92, 93, 94, 95, 96, 97, 98,
  99, 100, 101, 102, 103, 104, 105, 106, 107, 108, 109,
  110, 111, 112, 113, 114, 115, 116, 117, 118, 119, 120,
  121, 122, 123, 124, 125, 126, 127, 128, 129, 130, 131,
  132, 133, 134, 135, 136, 137, 138, 139, 140, 141, 142,
  143, 144, 145, 146, 147, 148, 149, 150, 151, 152, 153,
  154, 155, 156, 157, 158, 159, 160, 161, 162, 163, 164,
  165, 166, 167, 168, 169, 170, 171, 172, 173, 174, 175,
  176, 177, 178, 179, 180, 181, 182, 183, 184, 185, 186,
  187, 188, 189, 190, 191, 192, 193, 194, 195, 196, 197,
  198, 199, 200, 201, 202, 203, 204, 205, 206, 207, 208,
  209, 210, 211, 212, 213, 214, 215, 216, 217, 218, 219,
  220, 221, 222, 223, 224, 225, 226, 227, 228, 229, 230,
  231, 232, 233, 234, 235, 236, 237, 238, 239, 240, 241,
  242, 243, 244, 245, 246, 247, 248, 249, 250, 251, 252,
  253, 254, 255, 256, 257, 258, 259, 260, 261, 262, 263,
  264, 265, 266, 267, 268, 269, 270, 271, 272, 273, 274,
  275, 276, 277, 278, 279, 280, 281, 282, 283, 284, 285,
  286, 287, 288, 289, 290, 291, 292, 293, 294, 295, 296,
  297, 298, 299, 300, 301, 302, 303, 304, 305, 306, 307,
  308, 309, 310, 311, 312, 313, 314, 315, 316, 317, 318,
  319, 320, 321, 322, 323, 324, 325, 326, 327, 328, 329,
  330, 331, 332, 333, 334, 335, 336, 337, 338, 339, 340,
  341, 342, 343, 344, 345, 346, 347, 348, 349, 350, 351,
  352, 353, 354, 355, 356, 357, 358, 359, 360, 361, 362,
  363, 364, 365, 366, 367, 368, 369, 370, 371, 372, 373,
  374, 375, 376, 377, 378, 379, 380, 381, 382, 383, 384,
  385, 386, 387, 388, 389, 390, 391, 392, 393, 394, 395,
  396, 397, 398, 399, 400, 401, 402, 403, 404, 405, 406,
  407, 408, 409, 410, 411, 412, 413, 414, 415, 416, 417,
  418, 419, 420, 421, 422, 423, 424, 425, 426, 427, 428,
  429, 430, 431, 432, 433, 434, 435, 436, 437, 438, 439,
  440, 441, 442, 443, 444, 445, 446, 447, 448, 449, 450,
  451, 452, 453, 454, 455, 456, 457, 458, 459, 460, 461,
  462, 463, 464, 465, 466, 467, 468, 469, 470, 471, 472,
  473, 474, 475, 476, 477, 478, 479, 480, 481, 482, 483,
  484, 485, 486, 487, 488, 489, 490, 491, 492, 493, 494,
  495, 496, 497, 498, 499, 500, 501, 502, 503, 504, 505,
  506, 507, 508, 509, 510, 511, 512, 513, 514, 515, 516,
  517, 518, 519, 520, 521, 522, 523, 524, 525, 526, 527,
  528, 529, 530, 531, 532, 533, 534, 535, 536, 537, 538,
  539, 540, 541, 542, 543, 544, 545, 546, 547, 548, 549,
  550, 551, 552, 553, 554, 555, 556, 557, 558, 559, 560,
  561, 562, 563, 564, 565, 566, 567, 568, 569, 570, 571,
  572, 573, 574, 575, 576, 577, 578, 579, 580, 581, 582,
  583, 584, 585, 586, 587, 588, 589, 590, 591, 592, 593,
  594, 595, 596, 597, 598, 599, 600, 601, 602, 603, 604,
  605, 606, 607, 608, 609, 610, 611, 612, 613, 614, 615,
  616, 617, 618, 619, 620, 621, 622, 623, 624, 625, 626,
  627, 628, 629, 630, 631, 632, 633, 634, 635, 636, 637,
  638, 639, 640, 641, 642, 643, 644, 645, 646, 647, 648,
  649, 650, 651, 652, 653, 654, 655, 656, 657, 658, 659,
  660, 661, 662, 663, 664, 665, 666, 667, 668, 669, 670,
  671, 672, 673, 674, 675, 676, 677, 678, 679, 680, 681,
  682, 683, 684, 685, 686, 687, 688, 689, 690, 691, 692,
  693, 694, 695, 696, 697, 698, 699, 700, 701, 702, 703,
  704, 705, 706, 707, 708, 709, 710, 711, 712, 713, 714,
  715, 716, 717, 718, 719, 720, 721, 722, 723, 724, 725,
  726, 727, 728, 729, 730, 731, 732, 733, 734, 735, 736,
  737, 738, 739, 740, 741, 742, 743, 744, 745, 746, 747,
  748, 749, 750, 751, 752, 753, 754, 755, 756, 757, 758,
  759, 760, 761, 762, 763, 764, 765, 766, 767, 768, 769,
  770, 771, 772, 773, 774, 775, 776, 777, 778, 779, 780,
  781, 782, 783, 784, 785, 786, 787, 788, 789, 790, 791,
  792, 793, 794, 795, 796, 797, 798, 799, 800, 801, 802,
  803, 804, 805, 806, 807, 808, 809, 810, 811, 812, 813,
  814, 815, 816, 817, 818, 819, 820, 821, 822, 823, 824,
  825, 826, 827, 828, 829, 830, 831, 832, 833, 834, 835,
  836, 837, 838, 839, 840, 841, 842, 843, 844, 845, 846,
  847, 848, 849, 850, 851, 852, 853, 854, 855, 856, 857,
  858, 859, 860, 861, 862, 863, 864, 865, 866, 867, 868,
  869, 870, 871, 872, 873, 874, 875, 876, 877, 878, 879,
  880, 881, 882, 883, 884, 885, 886, 887, 888, 889, 890,
  891, 892, 893, 894, 895, 896, 897, 898, 899, 900, 901,
  902, 903, 904, 905, 906, 907, 908, 909, 910, 911, 912,
  913, 914, 915, 916, 917, 918, 919, 920, 921, 922, 923,
  924, 925, 926, 927, 928, 929, 930, 931, 932, 933, 934,
  935, 936, 937, 938, 939, 940, 941, 942, 943, 944, 945,
  946, 947, 948, 949, 950, 951, 952, 953, 954, 955, 956,
  957, 958, 959, 960, 961, 962, 963, 964, 965, 966, 967,
  968, 969, 970, 971, 972, 973, 974, 975, 976, 977, 978,
  979, 980, 981, 982, 983, 984, 985, 986, 987, 988, 989,
  990, 991, 992, 993, 994, 995, 996, 997, 998, 999, 1000,
  1001, 1002, 1003, 1004, 1005, 1006, 1007, 1008, 1009, 1010, 1011,
  1012, 1013, 1014, 1015, 1016, 1017, 1018, 1019, 1020, 1021, 1022,
  1023, 1024, 1025, 1026, 1027, 1028, 1029, 1030, 1031, 1032, 1033,
  1034, 1035, 1036, 1037, 1038, 1039, 1040, 1041, 1042, 1043, 1044,
  1045, 1046, 1047, 1048, 1049, 1050, 1051, 1052, 1053, 1054, 1055,
  1056, 1057, 1058, 1059, 1060, 1061, 1062, 1063, 1064, 1065, 1066,
  1067, 1068, 1069, 1070, 1071, 1072, 1073, 1074, 1075, 1076, 1077,
  1078, 1079, 1080, 1081, 1082, 1083, 1084, 1085, 1086, 1087, 1088,
  1089, 1090, 1091, 1092, 1093, 1094, 1095, 1096, 1097, 1098, 1099,
  1100, 1101, 1102, 1103, 1104, 1105, 1106, 1107, 1108, 1109, 1110,
  1111, 1112, 1113, 1114, 1115, 1116, 1117, 1118, 1119, 1120, 1121,
  1122, 1123, 1124, 1125, 1126, 1127, 1128, 1129, 1130, 1131, 1132,
  1133, 1134, 1135, 1136, 1137, 1138, 1139, 1140, 1141, 1142, 1143,
  1144, 1145, 1146, 1147, 1148, 1149, 1150, 1151, 1152, 1153, 1154,
  1155, 1156, 1157, 1158, 1159, 1160, 1161, 1162, 1163, 1164, 1165,
  1166, 1167, 1168, 1169, 1170, 1171, 1172, 1173, 1174, 1175, 1176,
  1177, 1178, 1179, 1180, 1181, 1182, 1183, 1184, 1185, 1186, 1187,
  1188, 1189, 1190, 1191, 1192, 1193, 1194, 1195, 1196, 1197, 1198,
  1199, 1200, 1201, 1202, 1203, 1204, 1205, 1206, 1207, 1208, 1209,
  1210, 1211, 1212, 1213, 1214, 1215, 1216, 1217, 1218, 1219, 1220,
  1221, 1222, 1223, 1224, 1225, 1226, 1227, 1228, 1229, 1230, 1231,
  1232, 1233, 1234, 1235, 1236, 1237, 1238, 1239, 1240, 1241, 1242,
  1243, 1244, 1245, 1246, 1247, 1248, 1249, 1250, 1251, 1252, 1253,
  1254, 1255, 1256, 1257, 1258, 1259, 1260, 1261, 1262, 1263, 1264,
  1265, 1266, 1267, 1268, 1269, 1270, 1271, 1272, 1273, 1274, 1275,
  1276, 1277, 1278, 1279, 1280, 1281, 1282, 1283, 1284, 1285, 1286,
  1287, 1288, 1289, 1290, 1291, 1292, 1293, 1294, 1295, 1296, 1297,
  1298, 1299, 1300, 1301, 1302, 1303, 1304, 1305, 1306, 1307, 1308,
  1309, 1310, 1311, 1312, 1313, 1314, 1315, 1316, 1317, 1318, 1319,
  1320, 1321, 1322, 1323, 1324, 1325, 1326, 1327, 1328, 1329, 1330,
  1331, 1332, 1333, 1334, 1335, 1336, 1337, 1338, 1339, 1340, 1341,
  1342, 1343, 1344, 1345, 1346, 1347, 1348, 1349, 1350, 1351, 1352,
  1353, 1354, 1355, 1356, 1357, 1358, 1359, 1360, 1361, 1362, 1363,
  1364, 1365, 1366, 1367, 1368, 1369, 1370, 1371, 1372, 1373, 1374,
  1375, 1376, 1377, 1378, 1379, 1380, 1381, 1382, 1383, 1384, 1385,
  1386, 1387, 1388, 1389, 1390, 1391, 1392, 1393, 1394, 1395, 1396,
  1397, 1398, 1399, 1400, 1401, 1402, 1403, 1404, 1405, 1406, 1407,
  1408, 1409, 1410, 1411, 1412, 1413, 1414, 1415, 1416, 1417, 1418,
  1419, 1420, 1421, 1422, 1423, 1424, 1425, 1426, 1427, 1428, 1429,
  1430, 1431, 1432, 1433, 1434, 1435, 1436, 1437, 1438, 1439, 1440,
  1441, 1442, 1443, 1444, 1445, 1446, 1447, 1448, 1449, 1450, 1451,
  1452, 1453, 1454, 1455, 1456, 1457, 1458, 1459, 1460, 1461, 1462,
  1463, 1464, 1465, 1466, 1467, 1468, 1469, 1470, 1471, 1472, 1473,
  1474, 1475, 1476, 1477, 1478, 1479, 1480, 1481, 1482, 1483, 1484,
  1485, 1486, 1487, 1488, 1489, 1490, 1491, 1492, 1493, 1494, 1495,
  1496, 1497, 1498, 1499, 1500, 1501, 1502, 1503, 1504, 1505, 1506,
  1507, 1508, 1509, 1510, 1511, 1512, 1513, 1514, 1515, 1516, 1517,
  1518, 1519, 1520, 1521, 1522, 1523, 1524, 1525, 1526, 1527, 1528,
  1529, 1530, 1531, 1532, 1533, 1534, 1535, 1536, 1537, 1538, 1539,
  1540, 1541, 1542, 1543, 1544, 1545, 1546, 1547, 1548, 1549, 1550,
  1551, 1552, 1553, 1554, 1555, 1556, 1557, 1558, 1559, 1560, 1561,
  1562, 1563, 1564, 1565, 1566, 1567, 1568, 1569, 1570, 1571, 1572,
  1573, 1574, 1575, 1576, 1577, 1578, 1579, 1580, 1581, 1582, 1583,
  1584, 1585, 1586, 1587, 1588, 1589, 1590, 1591, 1592, 1593, 1594,
  1595, 1596, 1597, 1598, 1599, 1600, 1601, 1602, 1603, 1604, 1605,
  1606, 1607, 1608, 1609, 1610, 1611, 1612, 1613, 1614, 1615, 1616,
  1617, 1618, 1619, 1620, 1621, 1622, 1623, 1624, 1625, 1626, 1627,
  1628, 1629, 1630, 1631, 1632, 1633, 1634, 1635, 1636, 1637, 1638,
  1639, 1640, 1641, 1642, 1643, 1644, 1645, 1646, 1647, 1648, 1649,
  1650, 1651, 1652, 1653, 1654, 1655, 1656, 1657, 1658, 1659, 1660,
  1661, 1662, 1663, 1664, 1665, 1666, 1667, 1668, 1669, 1670, 1671,
  1672, 1673, 1674, 1675, 1676, 1677, 1678, 1679, 1680, 1681, 1682,
  1683, 1684, 1685, 1686, 1687, 1688, 1689, 1690, 1691, 1692, 1693,
  1694, 1695, 1696, 1697, 1698, 1699, 1700, 1701, 1702, 1703, 1704,
  1705, 1706, 1707, 1708, 1709, 1710, 1711, 1712, 1713, 1714, 1715,
  1716, 1717, 1718, 1719, 1720, 1721, 1722, 1723, 1724, 1725, 1726,
  1727, 1728, 1729, 1730, 1731, 1732, 1733, 1734, 1735, 1736, 1737,
  1738, 1739, 1740, 1741, 1742, 1743, 1744, 1745, 1746, 1747, 1748,
  1749, 1750, 1751, 1752, 1753, 1754, 1755, 1756, 1757, 1758, 1759,
  1760, 1761, 1762, 1763, 1764, 1765, 1766, 1767, 1768, 1769, 1770,
  1771, 1772, 1773, 1774, 1775, 1776, 1777, 1778, 1779, 1780, 1781,
  1782, 1783, 1784, 1785, 1786, 1787, 1788, 1789, 1790, 1791, 1792,
  1793, 1794, 1795, 1796, 1797, 1798, 1799, 1800, 1801, 1802, 1803,
  1804, 1805, 1806, 1807, 1808, 1809, 1810, 1811, 1812, 1813, 1814,
  1815, 1816, 1817, 1818, 1819, 1820, 1821, 1822, 1823, 1824, 1825,
  1826, 1827, 1828, 1829, 1830, 1831, 1832, 1833, 1834, 1835, 1836,
  1837, 1838, 1839, 1840, 1841, 1842, 1843, 1844, 1845, 1846, 1847,
  1848, 1849, 1850, 1851, 1852, 1853, 1854, 1855, 1856, 1857, 1858,
  1859, 1860, 1861, 1862, 1863, 1864, 1865, 1866, 1867, 1868, 1869,
  1870, 1871, 1872, 1873, 1874, 1875, 1876, 1877, 1878, 1879, 1880,
  1881, 1882, 1883, 1884, 1885, 1886, 1887, 1888, 1889, 1890, 1891,
  1892, 1893, 1894, 1895, 1896, 1897, 1898, 1899, 1900, 1901, 1902,
  1903, 1904, 1905, 1906, 1907, 1908, 1909, 1910, 1911, 1912, 1913,
  1914, 1915, 1916, 1917, 1918, 1919, 1920, 1921, 1922, 1923, 1924,
  1925, 1926, 1927, 1928, 1929, 1930, 1931, 1932, 1933, 1934, 1935 ;

 sea_level_pressure =
  10168, 10164, 10158, 10152, 10146, 10138, 10130, 10124, 10118, 10112, 10101,
  10171, 10165, 10159, 10153, 10146, 10138, 10130, 10122, 10116, 10111, 10106,
  10172, 10166, 10161, 10154, 10147, 10139, 10131, 10123, 10115, 10109, 10107,
  10173, 10168, 10163, 10156, 10149, 10141, 10133, 10125, 10116, 10109, 10104,
  10176, 10171, 10166, 10159, 10152, 10145, 10137, 10129, 10121, 10112, 10103,
  10180, 10175, 10170, 10164, 10158, 10150, 10143, 10135, 10128, 10120, 10110,
  10184, 10180, 10175, 10168, 10162, 10156, 10150, 10143, 10135, 10129, 10122,
  10188, 10184, 10178, 10173, 10166, 10162, 10157, 10150, 10142, 10138, 10134,
  10193, 10187, 10182, 10177, 10171, 10167, 10162, 10155, 10150, 10146, 10143,
  10197, 10192, 10188, 10183, 10178, 10172, 10167, 10161, 10157, 10154, 10151,
  10202, 10197, 10194, 10190, 10185, 10179, 10173, 10168, 10164, 10161, 10158,
  10167, 10163, 10158, 10151, 10145, 10138, 10131, 10124, 10118, 10110, 10098,
  10170, 10164, 10159, 10152, 10146, 10138, 10130, 10123, 10117, 10111, 10106,
  10172, 10166, 10161, 10154, 10147, 10139, 10131, 10123, 10116, 10111, 10108,
  10174, 10169, 10163, 10156, 10148, 10141, 10133, 10125, 10117, 10110, 10105,
  10176, 10171, 10166, 10159, 10151, 10144, 10137, 10129, 10121, 10112, 10103,
  10179, 10175, 10169, 10163, 10157, 10150, 10143, 10135, 10127, 10118, 10109,
  10183, 10179, 10173, 10168, 10162, 10155, 10148, 10141, 10135, 10127, 10120,
  10187, 10183, 10178, 10172, 10166, 10160, 10154, 10148, 10142, 10136, 10132,
  10190, 10188, 10183, 10176, 10170, 10166, 10161, 10155, 10149, 10144, 10141,
  10195, 10193, 10188, 10182, 10175, 10171, 10166, 10161, 10156, 10152, 10149,
  10201, 10197, 10194, 10188, 10182, 10177, 10171, 10166, 10163, 10159, 10156,
  10166, 10163, 10157, 10150, 10145, 10139, 10131, 10125, 10119, 10109, 10095,
  10170, 10164, 10159, 10152, 10146, 10139, 10131, 10124, 10117, 10112, 10106,
  10172, 10166, 10160, 10154, 10147, 10139, 10131, 10124, 10117, 10112, 10109,
  10173, 10168, 10162, 10155, 10148, 10140, 10133, 10125, 10118, 10111, 10105,
  10175, 10170, 10164, 10157, 10151, 10144, 10136, 10128, 10120, 10112, 10103,
  10178, 10174, 10168, 10161, 10155, 10148, 10140, 10133, 10125, 10117, 10107,
  10182, 10177, 10172, 10166, 10160, 10153, 10145, 10138, 10132, 10125, 10117,
  10185, 10181, 10176, 10171, 10166, 10158, 10151, 10145, 10140, 10133, 10128,
  10189, 10185, 10182, 10176, 10170, 10163, 10157, 10152, 10147, 10142, 10137,
  10194, 10190, 10187, 10180, 10174, 10168, 10164, 10159, 10154, 10149, 10145,
  10199, 10196, 10192, 10186, 10179, 10174, 10170, 10166, 10161, 10157, 10153,
  10162, 10158, 10153, 10146, 10141, 10135, 10128, 10122, 10117, 10106, 10089,
  10166, 10160, 10154, 10148, 10141, 10134, 10128, 10121, 10114, 10109, 10102,
  10168, 10162, 10156, 10149, 10142, 10135, 10128, 10121, 10113, 10108, 10105,
  10169, 10164, 10157, 10151, 10144, 10137, 10129, 10121, 10113, 10107, 10100,
  10170, 10165, 10159, 10152, 10146, 10138, 10129, 10122, 10115, 10107, 10097,
  10174, 10169, 10163, 10156, 10149, 10142, 10134, 10126, 10119, 10112, 10101,
  10177, 10172, 10167, 10161, 10154, 10148, 10140, 10132, 10125, 10119, 10111,
  10181, 10176, 10171, 10166, 10160, 10154, 10147, 10139, 10133, 10128, 10122,
  10185, 10179, 10175, 10171, 10166, 10159, 10152, 10146, 10141, 10136, 10132,
  10190, 10185, 10181, 10177, 10171, 10165, 10159, 10154, 10149, 10144, 10140,
  10195, 10191, 10187, 10182, 10176, 10171, 10166, 10162, 10157, 10152, 10149 ;

 surface_snow_sickness =
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _ ;
}
